`timescale 1ns / 1ps

module tb_top();

    reg clk ,rst, btnU, btnD, echo, rx; 
    reg [3:0] sw;

    wire [3:0] fnd_com;
    wire [7:0] fnd_data;
    wire trig, tx;

    parameter us_10 = 10_000;
    parameter ms_1 = 1_000_000;

    Top u_top(
        .clk(clk),
        .rst(rst),
        .sw(sw),
        .sw_sub(),
        .btnU(btnU),
        .btnD(btnD),
        .btnL(),
        .btnR(),
        .echo(echo),
        .rx(rx),

        .fnd_com(fnd_com),
        .fnd_data(fnd_data),
        .trig(trig),
        .tx(tx),
        .led(),
        .sw_sub_led(),
        .watch_state_led(),

        .dht11_io()
    );

    always #5 clk = ~clk;

    initial begin
        #0; clk = 0; rst = 1; sw = 4'b0000; echo = 0; rx = 1; btnU = 0; btnD = 0;

        #20; rst = 0; sw = 4'b0100;
        #(10416 * 10);

        rx = 0;  // start
        #(10416 * 10);
        rx = 1;  // d0
        #(10416 * 10);
        rx = 1;  // d1
        #(10416 * 10);
        rx = 1;  // d2
        #(10416 * 10);
        rx = 0;  // d3
        #(10416 * 10);
        rx = 1;  // d4
        #(10416 * 10);
        rx = 0;  // d5
        #(10416 * 10);
        rx = 1;  // d6
        #(10416 * 10);
        rx = 0;  // d7
        #(10416 * 10);

        rx = 1;  // stop

        #50000;
        
        #25000;  //25us
        echo = 1'b1;
        #(1000*1000); // 1000ms
        echo = 1'b0;
        #25000;  //25us
        echo = 1'b1;
        #(1000*1000); // 1000ms
        echo = 1'b0;

        #ms_1;

        rx = 0;  // start
        #(10416 * 10);
        rx = 1;  // d0
        #(10416 * 10);
        rx = 1;  // d1
        #(10416 * 10);
        rx = 0;  // d2
        #(10416 * 10);
        rx = 0;  // d3
        #(10416 * 10);
        rx = 1;  // d4
        #(10416 * 10);
        rx = 0;  // d5
        #(10416 * 10);
        rx = 1;  // d6
        #(10416 * 10);
        rx = 0;  // d7
        #(10416 * 10);

        rx = 1;  // stop
        
        #ms_1;

        rx = 0;  // start
        #(10416 * 10);
        rx = 1;  // d0
        #(10416 * 10);
        rx = 1;  // d1
        #(10416 * 10);
        rx = 1;  // d2
        #(10416 * 10);
        rx = 0;  // d3
        #(10416 * 10);
        rx = 1;  // d4
        #(10416 * 10);
        rx = 0;  // d5
        #(10416 * 10);
        rx = 1;  // d6
        #(10416 * 10);
        rx = 0;  // d7
        #(10416 * 10);

        rx = 1;  // stop

        #ms_1;
        
        rx = 0;  // start
        #(10416 * 10);
        rx = 1;  // d0
        #(10416 * 10);
        rx = 1;  // d1
        #(10416 * 10);
        rx = 0;  // d2
        #(10416 * 10);
        rx = 0;  // d3
        #(10416 * 10);
        rx = 1;  // d4
        #(10416 * 10);
        rx = 1;  // d5
        #(10416 * 10);
        rx = 1;  // d6
        #(10416 * 10);
        rx = 1;  // d7
        #(10416 * 10);

        rx = 1;  // stop

        #ms_1;
        #50000;  //25us
        #25000;  //25us
        echo = 1'b1;
        #(1000*3000); // 1000ms
        echo = 1'b0;
        #25000;  //25us
        echo = 1'b1;
        #(1000*3000); // 1000ms
        echo = 1'b0;

        #ms_1;

        rx = 0;  // start
        #(10416 * 10);
        rx = 1;  // d0
        #(10416 * 10);
        rx = 1;  // d1
        #(10416 * 10);
        rx = 0;  // d2
        #(10416 * 10);
        rx = 0;  // d3
        #(10416 * 10);
        rx = 1;  // d4
        #(10416 * 10);
        rx = 0;  // d5
        #(10416 * 10);
        rx = 1;  // d6
        #(10416 * 10);
        rx = 0;  // d7
        #(10416 * 10);

        rx = 1;  // stop

        #ms_1;
        rx = 0;  // start
        #(10416 * 10);
        rx = 1;  // d0
        #(10416 * 10);
        rx = 1;  // d1
        #(10416 * 10);
        rx = 1;  // d2
        #(10416 * 10);
        rx = 0;  // d3
        #(10416 * 10);
        rx = 1;  // d4
        #(10416 * 10);
        rx = 0;  // d5
        #(10416 * 10);
        rx = 1;  // d6
        #(10416 * 10);
        rx = 0;  // d7
        #(10416 * 10);

        rx = 1;  // stop

        #50000;
        #25000;  //25us
        echo = 1'b1;
        #(1000*1000); // 1000ms
        echo = 1'b0;
        #25000;  //25us
        echo = 1'b1;
        #(1000*1000); // 1000ms
        echo = 1'b0;

        $stop;

    end
endmodule
